module decoder3_8(input [2:0]I,output [7:0]O);
assign O=1<<I;
endmodule
